// File name : lpsx_precalc.sv
// Version : 1.0
// Date : 1.03.2024
// URL : https://github.com/RomanVernin/streebog
// Author : Roman Vernin
`timescale 1ns/10ps
module lpsx_precalc #(
    parameter DATA_WIDTH = 512
)
(
    input   wire                            clk_i,
    input   wire                            rstn_i,
    input   wire                            valid_i,
    input   wire     [DATA_WIDTH-1:0]       lps_n_i,
    input   wire     [DATA_WIDTH-1:0]       lps_m_i,
    output  logic    [DATA_WIDTH-1:0]       lps_o,
    output  logic                           valid_o
);
logic [0:255] [63:0] T;
  
logic  [DATA_WIDTH-1:0] state_f;
logic [63:0][7:0]state;
logic [7:0] [DATA_WIDTH/8-1:0]  internal;
  
  //pre-calculation tables for pi, tau and L transformations
logic [0:255][63:0] T0 = {64'hd01f715b5c7ef8e6, 64'h16fa240980778325, 64'ha8a42e857ee049c8, 64'h6ac1068fa186465b,
      64'h6e417bd7a2e9320b, 64'h665c8167a437daab, 64'h7666681aa89617f6, 64'h4b959163700bdcf5,
      64'hf14be6b78df36248, 64'hc585bd689a625cff, 64'h9557d7fca67d82cb, 64'h89f0b969af6dd366,
      64'hb0833d48749f6c35, 64'ha1998c23b1ecbc7c, 64'h8d70c431ac02a736, 64'hd6dfbc2fd0a8b69e,
      64'h37aeb3e551fa198b, 64'h0b7d128a40b5cf9c, 64'h5a8f2008b5780cbc, 64'hedec882284e333e5,
      64'hd25fc177d3c7c2ce, 64'h5e0f5d50b61778ec, 64'h1d873683c0c24cb9, 64'had040bcbb45d208c,
      64'h2f89a0285b853c76, 64'h5732fff6791b8d58, 64'h3e9311439ef6ec3f, 64'hc9183a809fd3c00f,
      64'h83adf3f5260a01ee, 64'ha6791941f4e8ef10, 64'h103ae97d0ca1cd5d, 64'h2ce948121dee1b4a,
      64'h39738421dbf2bf53, 64'h093da2a6cf0cf5b4, 64'hcd9847d89cbcb45f, 64'hf9561c078b2d8ae8,
      64'h9c6a755a6971777f, 64'hbc1ebaa0712ef0c5, 64'h72e61542abf963a6, 64'h78bb5fde229eb12e,
      64'h14ba94250fceb90d, 64'h844d6697630e5282, 64'h98ea08026a1e032f, 64'hf06bbea144217f5c,
      64'hdb6263d11ccb377a, 64'h641c314b2b8ee083, 64'h320e96ab9b4770cf, 64'h1ee7deb986a96b85,
      64'he96cf57a878c47b5, 64'hfdd6615f8842feb8, 64'hc83862965601dd1b, 64'h2ea9f83e92572162,
      64'hf876441142ff97fc, 64'heb2c455608357d9d, 64'h5612a7e0b0c9904c, 64'h6c01cbfb2d500823,
      64'h4548a6a7fa037a2d, 64'habc4c6bf388b6ef4, 64'hbade77d4fdf8bebd, 64'h799b07c8eb4cac3a,
      64'h0c9d87e805b19cf0, 64'hcb588aac106afa27, 64'hea0c1d40c1e76089, 64'h2869354a1e816f1a,
      64'hff96d17307fbc490, 64'h9f0a9d602f1a5043, 64'h96373fc6e016a5f7, 64'h5292dab8b3a6e41c,
      64'h9b8ae0382c752413, 64'h4f15ec3b7364a8a5, 64'h3fb349555724f12b, 64'hc7c50d4415db66d7,
      64'h92b7429ee379d1a7, 64'hd37f99611a15dfda, 64'h231427c05e34a086, 64'ha439a96d7b51d538,
      64'hb403401077f01865, 64'hdda2aea5901d7902, 64'h0a5d4a9c8967d288, 64'hc265280adf660f93,
      64'h8bb0094520d4e94e, 64'h2a29856691385532, 64'h42a833c5bf072941, 64'h73c64d54622b7eb2,
      64'h07e095624504536c, 64'h8a905153e906f45a, 64'h6f6123c16b3b2f1f, 64'hc6e55552dc097bc3,
      64'h4468feb133d16739, 64'he211e7f0c7398829, 64'ha2f96419f7879b40, 64'h19074bdbc3ad38e9,
      64'hf4ebc3f9474e0b0c, 64'h43886bd376d53455, 64'hd8028beb5aa01046, 64'h51f23282f5cdc320,
      64'he7b1c2be0d84e16d, 64'h081dfab006dee8a0, 64'h3b33340d544b857b, 64'h7f5bcabc679ae242,
      64'h0edd37c48a08a6d8, 64'h81ed43d9a9b33bc6, 64'hb1a3655ebd4d7121, 64'h69a1eeb5e7ed6167,
      64'hf6ab73d5c8f73124, 64'h1a67a3e185c61fd5, 64'h2dc91004d43c065e, 64'h0240b02c8fb93a28,
      64'h90f7f2b26cc0eb8f, 64'h3cd3a16f114fd617, 64'haae49ea9f15973e0, 64'h06c0cd748cd64e78,
      64'hda423bc7d5192a6e, 64'hc345701c16b41287, 64'h6d2193ede4821537, 64'hfcf639494190e3ac,
      64'h7c3b228621f1c57e, 64'hfb16ac2b0494b0c0, 64'hbf7e529a3745d7f9, 64'h6881b6a32e3f7c73,
      64'hca78d2bad9b8e733, 64'hbbfe2fc2342aa3a9, 64'h0dbddffecc6381e4, 64'h70a6a56e2440598e,
      64'he4d12a844befc651, 64'h8c509c2765d0ba22, 64'hee8c6018c28814d9, 64'h17da7c1f49a59e31,
      64'h609c4c1328e194d3, 64'hb3e3d57232f44b09, 64'h91d7aaa4a512f69b, 64'h0ffd6fd243dabbcc,
      64'h50d26a943c1fde34, 64'h6be15e9968545b4f, 64'h94778fea6faf9fdf, 64'h2b09dd7058ea4826,
      64'h677cd9716de5c7bf, 64'h49d5214fffb2e6dd, 64'h0360e83a466b273c, 64'h1fc786af4f7b7691,
      64'ha0b9d435783ea168, 64'hd49f0c035f118cb6, 64'h01205816c9d21d14, 64'hac2453dd7d8f3d98,
      64'h545217cc3f70aa64, 64'h26b4028e9489c9c2, 64'hdec2469fd6765e3e, 64'h04807d58036f7450,
      64'he5f17292823ddb45, 64'hf30b569b024a5860, 64'h62dcfc3fa758aefb, 64'he84cad6c4e5e5aa1,
      64'hccb81fce556ea94b, 64'h53b282ae7a74f908, 64'h1b47fbf74c1402c1, 64'h368eebf39828049f,
      64'h7afbeff2ad278b06, 64'hbe5e0a8cfe97caed, 64'hcfd8f7f413058e77, 64'hf78b2bc301252c30,
      64'h4d555c17fcdd928d, 64'h5f2f05467fc565f8, 64'h24f4b2a21b30f3ea, 64'h860dd6bbecb768aa,
      64'h4c750401350f8f99, 64'h0000000000000000, 64'hecccd0344d312ef1, 64'hb5231806be220571,
      64'hc105c030990d28af, 64'h653c695de25cfd97, 64'h159acc33c61ca419, 64'hb89ec7f872418495,
      64'ha9847693b73254dc, 64'h58cf90243ac13694, 64'h59efc832f3132b80, 64'h5c4fed7c39ae42c4,
      64'h828dabe3efd81cfa, 64'hd13f294d95ace5f2, 64'h7d1b7a90e823d86a, 64'hb643f03cf849224d,
      64'h3df3f979d89dcb03, 64'h7426d836272f2dde, 64'hdfe21e891fa4432a, 64'h3a136c1b9d99986f,
      64'hfa36f43dcd46add4, 64'hc025982650df35bb, 64'h856d3e81aadc4f96, 64'hc4a5e57e53b041eb,
      64'h4708168b75ba4005, 64'haf44bbe73be41aa4, 64'h971767d029c4b8e3, 64'hb9be9feebb939981,
      64'h215497ecd18d9aae, 64'h316e7e91dd2c57f3, 64'hcef8afe2dad79363, 64'h3853dc371220a247,
      64'h35ee03c9de4323a3, 64'he6919aa8c456fc79, 64'he05157dc4880b201, 64'h7bdbb7e464f59612,
      64'h127a59518318f775, 64'h332ecebd52956ddb, 64'h8f30741d23bb9d1e, 64'hd922d3fd93720d52,
      64'h7746300c61440ae2, 64'h25d4eab4d2e2eefe, 64'h75068020eefd30ca, 64'h135a01474acaea61, 
      64'h304e268714fe4ae7, 64'ha519f17bb283c82c, 64'hdc82f6b359cf6416, 64'h5baf781e7caa11a8, 
      64'hb2c38d64fb26561d, 64'h34ce5bdf17913eb7, 64'h5d6fb56af07c5fd0, 64'h182713cd0a7f25fd,
      64'h9e2ac576e6c84d57, 64'h9aaab82ee5a73907, 64'ha3d93c0f3e558654, 64'h7e7b92aaae48ff56,
      64'h872d8ead256575be, 64'h41c8dbfff96c0e7d, 64'h99ca5014a3cc1e3b, 64'h40e883e930be1369,
      64'h1ca76e95091051ad, 64'h4e35b42dbab6b5b1, 64'h05a0254ecabd6944, 64'he1710fca8152af15,
      64'hf22b0e8dcb984574, 64'hb763a82a319b3f59, 64'h63fca4296e8ab3ef, 64'h9d4a2d4ca0a36a6b,
      64'he331bfe60eeb953d, 64'hd5bf541596c391a2, 64'hf5cb9bef8e9c1618, 64'h46284e9dbc685d11,
      64'h2074cffa185f87ba, 64'hbd3ee2b6b8fcedd1, 64'hae64e3f1f23607b0, 64'hfeb68965ce29d984,
      64'h55724fdaf6a2b770, 64'h29496d5cd753720e, 64'ha75941573d3af204, 64'h8e102c0bea69800a,
      64'h111ab16bc573d049, 64'hd7ffe439197aab8a, 64'hefac380e0b5a09cd, 64'h48f579593660fbc9,
      64'h22347fd697e6bd92, 64'h61bc1405e13389c7, 64'h4ab5c975b9d9c1e1, 64'h80cd1bcf606126d2,
      64'h7186fd78ed92449a, 64'h93971a882aabccb3, 64'h88d0e17f66bfce72, 64'h27945a985d5bd4d6
  };

logic [0:255][63:0] T1 = {64'hde553f8c05a811c8,64'h1906b59631b4f565,64'h436e70d6b1964ff7,64'h36d343cb8b1e9d85,
        64'h843dfacc858aab5a,64'hfdfc95c299bfc7f9,64'h0f634bdea1d51fa2,64'h6d458b3b76efb3cd,
        64'h85c3f77cf8593f80,64'h3c91315fbe737cb2,64'h2148b03366ace398,64'h18f8b8264c6761bf,  
        64'hc830c1c495c9fb0f,64'h981a76102086a0aa,64'haa16012142f35760,64'h35cc54060c763cf6,
        64'h42907d66cc45db2d,64'h8203d44b965af4bc,64'h3d6f3cefc3a0e868,64'hbc73ff69d292bda7,
        64'h8722ed0102e20a29,64'h8f8185e8cd34deb7,64'h9b0561dda7ee01d9,64'h5335a0193227fad6,
        64'hc9cecc74e81a6fd5,64'h54f5832e5c2431ea,64'h99e47ba05d553470,64'hf7bee756acd226ce,
        64'h384e05a5571816fd,64'hd1367452a47d0e6a,64'hf29fde1c386ad85b,64'h320c77316275f7ca,
        64'hd0c879e2d9ae9ab0,64'hdb7406c69110ef5d,64'h45505e51a2461011,64'hfc029872e46c5323,
        64'hfa3cb6f5f7bc0cc5,64'h031f17cd8768a173,64'hbd8df2d9af41297d,64'h9d3b4f5ab43e5e3f,
        64'h4071671b36feee84,64'h716207e7d3e3b83d,64'h48d20ff2f9283a1a,64'h27769eb4757cbc7e,
        64'h5c56ebc793f2e574,64'ha48b474f9ef5dc18,64'h52cbada94ff46e0c,64'h60c7da982d8199c6,
        64'h0e9d466edc068b78,64'h4eec2175eaf865fc,64'h550b8e9e21f7a530,64'h6b7ba5bc653fec2b,
        64'h5eb7f1ba6949d0dd,64'h57ea94e3db4c9099,64'hf640eae6d101b214,64'hdd4a284182c0b0bb,
        64'hff1d8fbf6304f250,64'hb8accb933bf9d7e8,64'he8867c478eb68c4d,64'h3f8e2692391bddc1,
        64'hcb2fd60912a15a7c,64'haec935dbab983d2f,64'hf55ffd2b56691367,64'h80e2ce366ce1c115,
        64'h179bf3f8edb27e1d,64'h01fe0db07dd394da,64'hda8a0b76ecc37b87,64'h44ae53e1df9584cb,
        64'hb310b4b77347a205,64'hdfab323c787b8512,64'h3b511268d070b78e,64'h65e6e3d2b9396753,
        64'h6864b271e2574d58,64'h259784c98fc789d7,64'h02e11a7dfabb35a9,64'h8841a6dfa337158b,
        64'h7ade78c39b5dcdd0,64'hb7cf804d9a2cc84a,64'h20b6bd831b7f7742,64'h75bd331d3a88d272,
        64'h418f6aab4b2d7a5e,64'hd9951cbb6babdaf4,64'hb6318dfde7ff5c90,64'h1f389b112264aa83,
        64'h492c024284fbaec0,64'he33a0363c608f9a0,64'h2688930408af28a4,64'hc7538a1a341ce4ad,
        64'h5da8e677ee2171ae,64'h8c9e92254a5c7fc4,64'h63d8cd55aae938b5,64'h29ebd8daa97a3706,
        64'h959827b37be88aa1,64'h1484e4356adadf6e,64'ha7945082199d7d6b,64'hbf6ce8a455fa1cd4,
        64'h9cc542eac9edcae5,64'h79c16f0e1c356ca3,64'h89bfab6fdee48151,64'hd4174d1830c5f0ff,
        64'h9258048415eb419d,64'h6139d72850520d1c,64'h6a85a80c18ec78f1,64'hcd11f88e0171059a,
        64'hcceff53e7ca29140,64'hd229639f2315af19,64'h90b91ef9ef507434,64'h5977d28d074a1be1,
        64'h311360fce51d56b9,64'hc093a92d5a1f2f91,64'h1a19a25bb6dc5416,64'heb996b8a09de2d3e,
        64'hfee3820f1ed7668a,64'hd7085ad5b7ad518c,64'h7fff41890fe53345,64'hec5948bd67dde602,
        64'h2fd5f65dbaaa68e0,64'ha5754affe32648c2,64'hf8ddac880d07396c,64'h6fa491468c548664,
        64'h0c7c5c1326bdbed1,64'h4a33158f03930fb3,64'h699abfc19f84d982,64'he4fa2054a80b329c,
        64'h6707f9af438252fa,64'h08a368e9cfd6d49e,64'h47b1442c58fd25b8,64'hbbb3dc5ebc91769b,
        64'h1665fe489061eac7,64'h33f27a811fa66310,64'h93a609346838d547,64'h30ed6d4c98cec263,
        64'h1dd9816cd8df9f2a,64'h94662a03063b1e7b,64'h83fdd9fbeb896066,64'h7b207573e68e590a,
        64'h5f49fc0a149a4407,64'h343259b671a5a82c,64'hfbc2bb458a6f981f,64'hc272b350a0a41a38,
        64'h3aaf1fd8ada32354,64'h6cbb868b0b3c2717,64'ha2b569c88d2583fe,64'hf180c9d1bf027928,
        64'haf37386bd64ba9f5,64'h12bacab2790a8088,64'h4c0d3b0810435055,64'hb2eeb9070e9436df,
        64'hc5b29067cea7d104,64'hdcb425f1ff132461,64'h4f122cc5972bf126,64'hac282fa651230886,
        64'he7e537992f6393ef,64'he61b3a2952b00735,64'h709c0a57ae302ce7,64'he02514ae416058d3,
        64'hc44c9dd7b37445de,64'h5a68c5408022ba92,64'h1c278cdca50c0bf0,64'h6e5a9cf6f18712be,
        64'h86dce0b17f319ef3,64'h2d34ec2040115d49,64'h4bcd183f7e409b69,64'h2815d56ad4a9a3dc,
        64'h24698979f2141d0d,64'h0000000000000000,64'h1ec696a15fb73e59,64'hd86b110b16784e2e,
        64'h8e7f8858b0e74a6d,64'h063e2e8713d05fe6,64'he2c40ed3bbdb6d7a,64'hb1f1aeca89fc97ac,
        64'he1db191e3cb3cc09,64'h6418ee62c4eaf389,64'hc6ad87aa49cf7077,64'hd6f65765ca7ec556,
        64'h9afb6c6dda3d9503,64'h7ce05644888d9236,64'h8d609f95378feb1e,64'h23a9aa4e9c17d631,
        64'h6226c0e5d73aac6f,64'h56149953a69f0443,64'heeb852c09d66d3ab,64'h2b0ac2a753c102af,
        64'h07c023376e03cb3c,64'h2ccae1903dc2c993,64'hd3d76e2f5ec63bc3,64'h9e2458973356ff4c,
        64'ha66a5d32644ee9b1,64'h0a427294356de137,64'h783f62be61e6f879,64'h1344c70204d91452,
        64'h5b96c8f0fdf12e48,64'ha90916ecc59bf613,64'hbe92e5142829880e,64'h727d102a548b194e,
        64'h1be7afebcb0fc0cc,64'h3e702b2244c8491b,64'hd5e940a84d166425,64'h66f9f41f3e51c620,
        64'habe80c913f20c3ba,64'hf07ec461c2d1edf2,64'hf361d3ac45b94c81,64'h0521394a94b8fe95,
        64'hadd622162cf09c5c,64'he97871f7f3651897,64'hf4a1f09b2bba87bd,64'h095d6559b2054044,
        64'h0bbc7f2448be75ed,64'h2af4cf172e129675,64'h157ae98517094bb4,64'h9fda55274e856b96,
        64'h914713499283e0ee,64'hb952c623462a4332,64'h74433ead475b46a8,64'h8b5eb112245fb4f8,
        64'ha34b6478f0f61724,64'h11a5dd7ffe6221fb,64'hc16da49d27ccbb4b,64'h76a224d0bde07301,
        64'h8aa0bca2598c2022,64'h4df336b86d90c48f,64'hea67663a740db9e4,64'hef465f70e0b54771,
        64'h39b008152acb8227,64'h7d1e5bf4f55e06ec,64'h105bd0cf83b1b521,64'h775c2960c033e7db,
        64'h7e014c397236a79f,64'h811cc386113255cf,64'heda7450d1a0e72d8,64'h5889df3d7a998f3b,
        64'h2e2bfbedc779fc3a,64'hce0eef438619a4e9,64'h372d4e7bf6cd095f,64'h04df34fae96b6a4f,
        64'hf923a13870d4adb6,64'ha1aa7e050a4d228d,64'ha8f71b5cb84862c9,64'hb52e9a306097fde3,
        64'h0d8251a35b6e2a0b,64'h2257a7fee1c442eb,64'h73831d9a29588d94,64'h51d4ba64c89ccf7f,
        64'h502ab7d4b54f5ba5,64'h97793dce8153bf08,64'he5042de4d5d8a646,64'h9687307efc802bd2,
        64'ha05473b5779eb657,64'hb4d097801d446939,64'hcff0e2f3fbca3033,64'hc38cbee0dd778ee2,
        64'h464f499c252eb162,64'hcad1dbb96f72cea6,64'hba4dd1eec142e241,64'hb00fa37af42f0376
        };

logic [0:255][63:0] T2 = {64'hcce4cd3aa968b245, 64'h089d5484e80b7faf, 64'h638246c1b3548304, 64'hd2fe0ec8c2355492,
        64'ha7fbdf7ff2374eee, 64'h4df1600c92337a16, 64'h84e503ea523b12fb, 64'h0790bbfd53ab0c4a,
        64'h198a780f38f6ea9d, 64'h2ab30c8f55ec48cb, 64'he0f7fed6b2c49db5, 64'hb6ecf3f422cadbdc,
        64'h409c9a541358df11, 64'hd3ce8a56dfde3fe3, 64'hc3e9224312c8c1a0, 64'h0d6dfa58816ba507,
        64'hddf3e1b179952777, 64'h04c02a42748bb1d9, 64'h94c2abff9f2decb8, 64'h4f91752da8f8acf4,
        64'h78682befb169bf7b, 64'he1c77a48af2ff6c4, 64'h0c5d7ec69c80ce76, 64'h4cc1e4928fd81167,
        64'hfeed3d24d9997b62, 64'h518bb6dfc3a54a23, 64'h6dbf2d26151f9b90, 64'hb5bc624b05ea664f,
        64'he86aaa525acfe21a, 64'h4801ced0fb53a0be, 64'hc91463e6c00868ed, 64'h1027a815cd16fe43,
        64'hf67069a0319204cd, 64'hb04ccc976c8abce7, 64'hc0b9b3fc35e87c33, 64'hf380c77c58f2de65,
        64'h50bb3241de4e2152, 64'hdf93f490435ef195, 64'hf1e0d25d62390887, 64'haf668bfb1a3c3141,
        64'hbc11b251f00a7291, 64'h73a5eed47e427d47, 64'h25bee3f6ee4c3b2e, 64'h43cc0beb34786282,
        64'hc824e778dde3039c, 64'hf97d86d98a327728, 64'hf2b043e24519b514, 64'he297ebf7880f4b57,
        64'h3a94a49a98fab688, 64'h868516cb68f0c419, 64'heffa11af0964ee50, 64'ha4ab4ec0d517f37d,
        64'ha9c6b498547c567a, 64'h8e18424f80fbbbb6, 64'h0bcdc53bcf2bc23c, 64'h137739aaea3643d0,
        64'h2c1333ec1bac2ff0, 64'h8d48d3f0a7db0625, 64'h1e1ac3f26b5de6d7, 64'hf520f81f16b2b95e,
        64'h9f0f6ec450062e84, 64'h0130849e1deb6b71, 64'hd45e31ab8c7533a9, 64'h652279a2fd14e43f,
        64'h3209f01e70f1c927, 64'hbe71a770cac1a473, 64'h0e3d6be7a64b1894, 64'h7ec8148cff29d840,
        64'hcb7476c7fac3be0f, 64'h72956a4a63a91636, 64'h37f95ec21991138f, 64'h9e3fea5a4ded45f5,
        64'h7b38ba50964902e8, 64'h222e580bbde73764, 64'h61e253e0899f55e6, 64'hfc8d2805e352ad80,
        64'h35994be3235ac56d, 64'h09add01af5e014de, 64'h5e8659a6780539c6, 64'hb17c48097161d796,
        64'h026015213acbd6e2, 64'hd1ae9f77e515e901, 64'hb7dc776a3f21b0ad, 64'haba6a1b96eb78098,
        64'h9bcf4486248d9f5d, 64'h582666c536455efd, 64'hfdbdac9bfeb9c6f1, 64'hc47999be4163cdea,
        64'h765540081722a7ef, 64'h3e548ed8ec710751, 64'h3d041f67cb51bac2, 64'h7958af71ac82d40a,
        64'h36c9da5c047a78fe, 64'hed9a048e33af38b2, 64'h26ee7249c96c86bd, 64'h900281bdeba65d61,
        64'h11172c8bd0fd9532, 64'hea0abf73600434f8, 64'h42fc8f75299309f3, 64'h34a9cf7d3eb1ae1c,
        64'h2b838811480723ba, 64'h5ce64c8742ceef24, 64'h1adae9b01fd6570e, 64'h3c349bf9d6bad1b3,
        64'h82453c891c7b75c0, 64'h97923a40b80d512b, 64'h4a61dbf1c198765c, 64'hb48ce6d518010d3e,
        64'hcfb45c858e480fd6, 64'hd933cbf30d1e96ae, 64'hd70ea014ab558e3a, 64'hc189376228031742,
        64'h9262949cd16d8b83, 64'heb3a3bed7def5f89, 64'h49314a4ee6b8cbcf, 64'hdcc3652f647e4c06,
        64'hda635a4c2a3e2b3d, 64'h470c21a940f3d35b, 64'h315961a157d174b4, 64'h6672e81dda3459ac,
        64'h5b76f77a1165e36e, 64'h445cb01667d36ec8, 64'hc5491d205c88a69b, 64'h456c34887a3805b9,
        64'hffddb9bac4721013, 64'h99af51a71e4649bf, 64'ha15be01cbc7729d5, 64'h52db2760e485f7b0,
        64'h8c78576eba306d54, 64'hae560f6507d75a30, 64'h95f22f6182c687c9, 64'h71c5fbf54489aba5,
        64'hca44f259e728d57e, 64'h88b87d2ccebbdc8d, 64'hbab18d32be4a15aa, 64'h8be8ec93e99b611e,
        64'h17b713e89ebdf209, 64'hb31c5d284baa0174, 64'heeca9531148f8521, 64'hb8d198138481c348,
        64'h8988f9b2d350b7fc, 64'hb9e11c8d996aa839, 64'h5a4673e40c8e881f, 64'h1687977683569978,
        64'hbf4123eed72acf02, 64'h4ea1f1b3b513c785, 64'he767452be16f91ff, 64'h7505d1b730021a7c,
        64'ha59bca5ec8fc980c, 64'had069eda20f7e7a3, 64'h38f4b1bba231606a, 64'h60d2d77e94743e97,
        64'h9affc0183966f42c, 64'h248e6768f3a7505f, 64'hcdd449a4b483d934, 64'h87b59255751baf68,
        64'h1bea6d2e023d3c7f, 64'h6b1f12455b5ffcab, 64'h743555292de9710d, 64'hd8034f6d10f5fddf,
        64'hc6198c9f7ba81b08, 64'hbb8109aca3a17edb, 64'hfa2d1766ad12cabb, 64'hc729080166437079,
        64'h9c5fff7b77269317, 64'h0000000000000000, 64'h15d706c9a47624eb, 64'h6fdf38072fd44d72,
        64'h5fb6dd3865ee52b7, 64'ha33bf53d86bcff37, 64'he657c1b5fc84fa8e, 64'haa962527735cebe9,
        64'h39c43525bfda0b1b, 64'h204e4d2a872ce186, 64'h7a083ece8ba26999, 64'h554b9c9db72efbfa,
        64'hb22cd9b656416a05, 64'h96a2bedea5e63a5a, 64'h802529a826b0a322, 64'h8115ad363b5bc853,
        64'h8375b81701901eb1, 64'h3069e53f4a3a1fc5, 64'hbd2136cfede119e0, 64'h18bafc91251d81ec,
        64'h1d4a524d4c7d5b44, 64'h05f0aedc6960daa8, 64'h29e39d3072ccf558, 64'h70f57f6b5962c0d4,
        64'h989fd53903ad22ce, 64'hf84d024797d91c59, 64'h547b1803aac5908b, 64'hf0d056c37fd263f6,
        64'hd56eb535919e58d8, 64'h1c7ad6d351963035, 64'h2e7326cd2167f912, 64'hac361a443d1c8cd2,
        64'h697f076461942a49, 64'h4b515f6fdc731d2d, 64'h8ad8680df4700a6f, 64'h41ac1eca0eb3b460,
        64'h7d988533d80965d3, 64'ha8f6300649973d0b, 64'h7765c4960ac9cc9e, 64'h7ca801adc5e20ea2,
        64'hdea3700e5eb59ae4, 64'ha06b6482a19c42a4, 64'h6a2f96db46b497da, 64'h27def6d7d487edcc,
        64'h463ca5375d18b82a, 64'ha6cb5be1efdc259f, 64'h53eba3fef96e9cc1, 64'hce84d81b93a364a7,
        64'hf4107c810b59d22f, 64'h333974806d1aa256, 64'h0f0def79bba073e5, 64'h231edc95a00c5c15,
        64'he437d494c64f2c6c, 64'h91320523f64d3610, 64'h67426c83c7df32dd, 64'h6eefbc99323f2603,
        64'h9d6f7be56acdf866, 64'h5916e25b2bae358c, 64'h7ff89012e2c2b331, 64'h035091bf2720bd93,
        64'h561b0d22900e4669, 64'h28d319ae6f279e29, 64'h2f43a2533c8c9263, 64'hd09e1be9f8fe8270,
        64'hf740ed3e2c796fbc, 64'hdb53ded237d5404c, 64'h62b2c25faebfe875, 64'h0afd41a5d2c0a94d,
        64'h6412fd3ce0ff8f4e, 64'he3a76f6995e42026, 64'h6c8fa9b808f4f0e1, 64'hc2d9a6dd0f23aad1,
        64'h8f28c6d19d10d0c7, 64'h85d587744fd0798a, 64'ha20b71a39b579446, 64'h684f83fa7c7f4138,
        64'he507500adba4471d, 64'h3f640a46f19a6c20, 64'h1247bd34f7dd28a1, 64'h2d23b77206474481,
        64'h93521002cc86e0f2, 64'h572b89bc8de52d18, 64'hfb1d93f8b0f9a1ca, 64'he95a2ecc4724896b,
        64'h3ba420048511ddf9, 64'hd63e248ab6bee54b, 64'h5dd6c8195f258455, 64'h06a03f634e40673b,
        64'h1f2a476c76b68da6, 64'h217ec9b49ac78af7, 64'hecaa80102e4453c3, 64'h14e78257b99d4f9a
        };

logic [0:255][63:0] T3 = {64'h20329b2cc87bba05, 64'h4f5eb6f86546a531, 64'hd4f44775f751b6b1, 64'h8266a47b850dfa8b,
        64'hbb986aa15a6ca985, 64'hc979eb08f9ae0f99, 64'h2da6f447a2375ea1, 64'h1e74275dcd7d8576,
        64'hbc20180a800bc5f8, 64'hb4a2f701b2dc65be, 64'he726946f981b6d66, 64'h48e6c453bf21c94c,
        64'h42cad9930f0a4195, 64'hefa47b64aacccd20, 64'h71180a8960409a42, 64'h8bb3329bf6a44e0c,
        64'hd34c35de2d36dacc, 64'ha92f5b7cbc23dc96, 64'hb31a85aa68bb09c3, 64'h13e04836a73161d2,
        64'hb24dfc4129c51d02, 64'h8ae44b70b7da5acd, 64'he671ed84d96579a7, 64'ha4bb3417d66f3832,
        64'h4572ab38d56d2de8, 64'hb1b47761ea47215c, 64'he81c09cf70aba15d, 64'hffbdb872ce7f90ac, 
        64'ha8782297fd5dc857, 64'h0d946f6b6a4ce4a4, 64'he4df1f4f5b995138, 64'h9ebc71edca8c5762,
        64'h0a2c1dc0b02b88d9, 64'h3b503c115d9d7b91, 64'hc64376a8111ec3a2, 64'hcec199a323c963e4,
        64'hdc76a87ec58616f7, 64'h09d596e073a9b487, 64'h14583a9d7d560daf, 64'hf4c6dc593f2a0cb4,
        64'hdd21d19584f80236, 64'h4a4836983ddde1d3, 64'he58866a41ae745f9, 64'hf591a5b27e541875,
        64'h891dc05074586693, 64'h5b068c651810a89e, 64'ha30346bc0c08544f, 64'h3dbf3751c684032d,
        64'h2a1e86ec785032dc, 64'hf73f5779fca830ea, 64'hb60c05ca30204d21, 64'h0cc316802b32f065,
        64'h8770241bdd96be69, 64'hb861e18199ee95db, 64'hf805cad91418fcd1, 64'h29e70dccbbd20e82,
        64'hc7140f435060d763, 64'h0f3a9da0e8b0cc3b, 64'ha2543f574d76408e, 64'hbd7761e1c175d139,
        64'h4b1f4f737ca3f512, 64'h6dc2df1f2fc137ab, 64'hf1d05c3967b14856, 64'ha742bf3715ed046c,
        64'h654030141d1697ed, 64'h07b872abda676c7d, 64'h3ce84eba87fa17ec, 64'hc1fb0403cb79afdf,
        64'h3e46bc7105063f73, 64'h278ae987121cd678, 64'ha1adb4778ef47cd0, 64'h26dd906c5362c2b9,
        64'h05168060589b44e2, 64'hfbfc41f9d79ac08f, 64'h0e6de44ba9ced8fa, 64'h9feb08068bf243a3,
        64'h7b341749d06b129b, 64'h229c69e74a87929a, 64'he09ee6c4427c011b, 64'h5692e30e725c4c3a,
        64'hda99a33e5e9f6e4b, 64'h353dd85af453a36b, 64'h25241b4c90e0fee7, 64'h5de987258309d022,
        64'he230140fc0802984, 64'h93281e86a0c0b3c6, 64'hf229d719a4337408, 64'h6f6c2dd4ad3d1f34,
        64'h8ea5b2fbae3f0aee, 64'h8331dd90c473ee4a, 64'h346aa1b1b52db7aa, 64'hdf8f235e06042aa9,
        64'hcc6f6b68a1354b7b, 64'h6c95a6f46ebf236a, 64'h52d31a856bb91c19, 64'h1a35ded6d498d555,
        64'hf37eaef2e54d60c9, 64'h72e181a9a3c2a61c, 64'h98537aad51952fde, 64'h16f6c856ffaa2530,
        64'hd960281e9d1d5215, 64'h3a0745fa1ce36f50, 64'h0b7b642bf1559c18, 64'h59a87eae9aec8001,
        64'h5e100c05408bec7c, 64'h0441f98b19e55023, 64'hd70dcc5534d38aef, 64'h927f676de1bea707,
        64'h9769e70db925e3e5, 64'h7a636ea29115065a, 64'h468b201816ef11b6, 64'hab81a9b73edff409,
        64'hc0ac7de88a07bb1e, 64'h1f235eb68c0391b7, 64'h6056b074458dd30f, 64'hbe8eeac102f7ed67,
        64'hcd381283e04b5fba, 64'h5cbefecec277c4e3, 64'hd21b4c356c48ce0d, 64'h1019c31664b35d8c,
        64'h247362a7d19eea26, 64'hebe582efb3299d03, 64'h02aef2cb82fc289f, 64'h86275df09ce8aaa8,
        64'h28b07427faac1a43, 64'h38a9b7319e1f47cf, 64'hc82e92e3b8d01b58, 64'h06ef0b409b1978bc,
        64'h62f842bfc771fb90, 64'h9904034610eb3b1f, 64'hded85ab5477a3e68, 64'h90d195a663428f98,
        64'h5384636e2ac708d8, 64'hcbd719c37b522706, 64'hae9729d76644b0eb, 64'h7c8c65e20a0c7ee6,
        64'h80c856b007f1d214, 64'h8c0b40302cc32271, 64'hdbcedad51fe17a8a, 64'h740e8ae938dbdea0,
        64'ha615c6dc549310ad, 64'h19cc55f6171ae90b, 64'h49b1bdb8fe5fdd8d, 64'hed0a89af2830e5bf,
        64'h6a7aadb4f5a65bd6, 64'h7e22972988f05679, 64'hf952b3325566e810, 64'h39fecedadf61530e,
        64'h6101c99f04f3c7ce, 64'h2e5f7f6761b562ff, 64'hf08725d226cf5c97, 64'h63af3b54860fef51,
        64'h8ff2cb10ef411e2f, 64'h884ab9bb35267252, 64'h4df04433e7ba8dae, 64'h9afd8866d3690741,
        64'h66b9bb34de94abb3, 64'h9baaf18d92171380, 64'h543c11c5f0a064a5, 64'h17a1b1bdbed431f1,
        64'hb5f58eeaf3a2717f, 64'hc355f6c849858740, 64'hec5df044694ef17e, 64'hd83751f5dc6346d4,
        64'hfc4433520dfdacf2, 64'h0000000000000000, 64'h5a51f58e596ebc5f, 64'h3285aaf12e34cf16,
        64'h8d5c39db6dbd36b0, 64'h12b731dde64f7513, 64'h94906c2d7aa7dfbb, 64'h302b583aacc8e789,
        64'h9d45facd090e6b3c, 64'h2165e2c78905aec4, 64'h68d45f7f775a7349, 64'h189b2c1d5664fdca,
        64'he1c99f2f030215da, 64'h6983269436246788, 64'h8489af3b1e148237, 64'he94b702431d5b59c,
        64'h33d2d31a6f4adbd7, 64'hbfd9932a4389f9a6, 64'hb0e30e8aab39359d, 64'hd1e2c715afcaf253,
        64'h150f43763c28196e, 64'hc4ed846393e2eb3d, 64'h03f98b20c3823c5e, 64'hfd134ab94c83b833,
        64'h556b682eb1de7064, 64'h36c4537a37d19f35, 64'h7559f30279a5ca61, 64'h799ae58252973a04,
        64'h9c12832648707ffd, 64'h78cd9c6913e92ec5, 64'h1d8dac7d0effb928, 64'h439da0784e745554,
        64'h413352b3cc887dcb, 64'hbacf134a1b12bd44, 64'h114ebafd25cd494d, 64'h2f08068c20cb763e,
        64'h76a07822ba27f63f, 64'heab2fb04f25789c2, 64'he3676de481fe3d45, 64'h1b62a73d95e6c194,
        64'h641749ff5c68832c, 64'ha5ec4dfc97112cf3, 64'hf6682e92bdd6242b, 64'h3f11c59a44782bb2,
        64'h317c21d1edb6f348, 64'hd65ab5be75ad9e2e, 64'h6b2dd45fb4d84f17, 64'hfaab381296e4d44e,
        64'hd0b5befeeeb4e692, 64'h0882ef0b32d7a046, 64'h512a91a5a83b2047, 64'h963e9ee6f85bf724,
        64'h4e09cf132438b1f0, 64'h77f701c9fb59e2fe, 64'h7ddb1c094b726a27, 64'h5f4775ee01f5f8bd,
        64'h9186ec4d223c9b59, 64'hfeeac1998f01846d, 64'hac39db1ce4b89874, 64'hb75b7c21715e59e0,
        64'hafc0503c273aa42a, 64'h6e3b543fec430bf5, 64'h704f7362213e8e83, 64'h58ff0745db9294c0,
        64'h67eec2df9feabf72, 64'ha0facd9ccf8a6811, 64'hb936986ad890811a, 64'h95c715c63bd9cb7a,
        64'hca8060283a2c33c7, 64'h507de84ee9453486, 64'h85ded6d05f6a96f6, 64'h1cdad5964f81ade9,
        64'hd5a33e9eb62fa270, 64'h40642b588df6690a, 64'h7f75eec2c98e42b8, 64'h2cf18dace3494a60,
        64'h23cb100c0bf9865b, 64'heef3028febb2d9e1, 64'h4425d2d394133929, 64'haad6d05c7fa1e0c8,
        64'had6ea2f7a5c68cb5, 64'hc2028f2308fb9381, 64'h819f2f5b468fc6d5, 64'hc5bafd88d29cfffc,
        64'h47dc59f357910577, 64'h2b49ff07392e261d, 64'h57c59ae5332258fb, 64'h73b6f842e2bcb2dd,
        64'hcf96e04862b77725, 64'h4ca73dd8a6c4996f, 64'h015779eb417e14c1, 64'h37932a9176af8bf4
        };
logic [0:255][63:0] T4 = {64'h190a2c9b249df23e, 64'h2f62f8b62263e1e9, 64'h7a7f754740993655, 64'h330b7ba4d5564d9f,
        64'h4c17a16a46672582, 64'hb22f08eb7d05f5b8, 64'h535f47f40bc148cc, 64'h3aec5d27d4883037,
        64'h10ed0a1825438f96, 64'h516101f72c233d17, 64'h13cc6f949fd04eae, 64'h739853c441474bfd,
        64'h653793d90d3f5b1b, 64'h5240647b96b0fc2f, 64'h0c84890ad27623e0, 64'hd7189b32703aaea3,
        64'h2685de3523bd9c41, 64'h99317c5b11bffefa, 64'h0d9baa854f079703, 64'h70b93648fbd48ac5,
        64'ha80441fce30bc6be, 64'h7287704bdc36ff1e, 64'hb65384ed33dc1f13, 64'hd36417343ee34408,
        64'h39cd38ab6e1bf10f, 64'h5ab861770a1f3564, 64'h0ebacf09f594563b, 64'hd04572b884708530,
        64'h3cae9722bdb3af47, 64'h4a556b6f2f5cbaf2, 64'he1704f1f76c4bd74, 64'h5ec4ed7144c6dfcf,
        64'h16afc01d4c7810e6, 64'h283f113cd629ca7a, 64'haf59a8761741ed2d, 64'heed5a3991e215fac, 
        64'h3bf37ea849f984d4, 64'he413e096a56ce33c, 64'h2c439d3a98f020d1, 64'h637559dc6404c46b,
        64'h9e6c95d1e5f5d569, 64'h24bb9836045fe99a, 64'h44efa466dac8ecc9, 64'hc6eab2a5c80895d6,
        64'h803b50c035220cc4, 64'h0321658cba93c138, 64'h8f9ebc465dc7ee1c, 64'hd15a5137190131d3,
        64'h0fa5ec8668e5e2d8, 64'h91c979578d1037b1, 64'h0642ca05693b9f70, 64'hefca80168350eb4f,
        64'h38d21b24f36a45ec, 64'hbeab81e1af73d658, 64'h8cbfd9cae7542f24, 64'hfd19cc0d81f11102,
        64'h0ac6430fbb4dbc90, 64'h1d76a09d6a441895, 64'h2a01573ff1cbbfa1, 64'hb572e161894fde2b,
        64'h8124734fa853b827, 64'h614b1fdf43e6b1b0, 64'h68ac395c4238cc18, 64'h21d837bfd7f7b7d2,
        64'h20c714304a860331, 64'h5cfaab726324aa14, 64'h74c5ba4eb50d606e, 64'hf3a3030474654739,
        64'h23e671bcf015c209, 64'h45f087e947b9582a, 64'hd8bd77b418df4c7b, 64'he06f6c90ebb50997,
        64'h0bd96080263c0873, 64'h7e03f9410e40dcfe, 64'hb8e94be4c6484928, 64'hfb5b0608e8ca8e72,
        64'h1a2b49179e0e3306, 64'h4e29e76961855059, 64'h4f36c4e6fcf4e4ba, 64'h49740ee395cf7bca,
        64'hc2963ea386d17f7d, 64'h90d65ad810618352, 64'h12d34c1b02a1fa4d, 64'hfa44258775bb3a91,
        64'h18150f14b9ec46dd, 64'h1491861e6b9a653d, 64'h9a1019d7ab2c3fc2, 64'h3668d42d06fe13d7,
        64'hdcc1fbb25606a6d0, 64'h969490dd795a1c22, 64'h3549b1a1bc6dd2ef, 64'hc94f5e23a0ed770e,
        64'hb9f6686b5b39fdcb, 64'hc4d4f4a6efeae00d, 64'he732851a1fff2204, 64'h94aad6de5eb869f9,
        64'h3f8ff2ae07206e7f, 64'hfe38a9813b62d03a, 64'ha7a1ad7a8bee2466, 64'h7b6056c8dde882b6,
        64'h302a1e286fc58ca7, 64'h8da0fa457a259bc7, 64'hb3302b64e074415b, 64'h5402ae7eff8b635f,
        64'h08f8050c9cafc94b, 64'hae468bf98a3059ce, 64'h88c355cca98dc58f, 64'hb10e6d67c7963480,
        64'hbad70de7e1aa3cf3, 64'hbfb4a26e320262bb, 64'hcb711820870f02d5, 64'hce12b7a954a75c9d,
        64'h563ce87dd8691684, 64'h9f73b65e7884618a, 64'h2b1e74b06cba0b42, 64'h47cec1ea605b2df1,
        64'h1c698312f735ac76, 64'h5fdbcefed9b76b2c, 64'h831a354c8fb1cdfc, 64'h820516c312c0791f,
        64'hb74ca762aeadabf0, 64'hfc06ef821c80a5e1, 64'h5723cbf24518a267, 64'h9d4df05d5f661451,
        64'h588627742dfd40bf, 64'hda8331b73f3d39a0, 64'h17b0e392d109a405, 64'hf965400bcf28fba9,
        64'h7c3dbf4229a2a925, 64'h023e460327e275db, 64'h6cd0b55a0ce126b3, 64'he62da695828e96e7,
        64'h42ad6e63b3f373b9, 64'he50cc319381d57df, 64'hc5cbd729729b54ee, 64'h46d1e265fd2a9912,
        64'h6428b056904eeff8, 64'h8be23040131e04b7, 64'h6709d5da2add2ec0, 64'h075de98af44a2b93,
        64'h8447dcc67bfbe66f, 64'h6616f655b7ac9a23, 64'hd607b8bded4b1a40, 64'h0563af89d3a85e48,
        64'h3db1b4ad20c21ba4, 64'h11f22997b8323b75, 64'h292032b34b587e99, 64'h7f1cdace9331681d,
        64'h8e819fc9c0b65aff, 64'ha1e3677fe2d5bb16, 64'hcd33d225ee349da5, 64'hd9a2543b85aef898,
        64'h795e10cbfa0af76d, 64'h25a4bbb9992e5d79, 64'h78413344677b438e, 64'hf0826688cef68601,
        64'hd27b34bba392f0eb, 64'h551d8df162fad7bc, 64'h1e57c511d0d7d9ad, 64'hdeffbdb171e4d30b,
        64'hf4feea8e802f6caa, 64'ha480c8f6317de55e, 64'ha0fc44f07fa40ff5, 64'h95b5f551c3c9dd1a,
        64'h22f952336d6476ea, 64'h0000000000000000, 64'ha6be8ef5169f9085, 64'hcc2cf1aa73452946,
        64'h2e7ddb39bf12550a, 64'hd526dd3157d8db78, 64'h486b2d6c08becf29, 64'h9b0f3a58365d8b21,
        64'hac78cdfaadd22c15, 64'hbc95c7e28891a383, 64'h6a927f5f65dab9c3, 64'hc3891d2c1ba0cb9e,
        64'heaa92f9f50f8b507, 64'hcf0d9426c9d6e87e, 64'hca6e3baf1a7eb636, 64'hab25247059980786,
        64'h69b31ad3df4978fb, 64'he2512a93cc577c4c, 64'hff278a0ea61364d9, 64'h71a615c766a53e26,
        64'h89dc764334fc716c, 64'hf87a638452594f4a, 64'hf2bc208be914f3da, 64'h8766b94ac1682757,
        64'hbbc82e687cdb8810, 64'h626a7a53f9757088, 64'ha2c202f358467a2e, 64'h4d0882e5db169161,
        64'h09e7268301de7da8, 64'he897699c771ac0dc, 64'hc8507dac3d9cc3ed, 64'hc0a878a0a1330aa6,
        64'h978bb352e42ba8c1, 64'he9884a13ea6b743f, 64'h279afdbabecc28a2, 64'h047c8c064ed9eaab,
        64'h507e2278b15289f4, 64'h599904fbb08cf45c, 64'hbd8ae46d15e01760, 64'h31353da7f2b43844,
        64'h8558ff49e68a528c, 64'h76fbfc4d92ef15b5, 64'h3456922e211c660c, 64'h86799ac55c1993b4,
        64'h3e90d1219a51da9c, 64'h2d5cbeb505819432, 64'h982e5fd48cce4a19, 64'hdb9c1238a24c8d43,
        64'hd439febecaa96f9b, 64'h418c0bef0960b281, 64'h158ea591f6ebd1de, 64'h1f48e69e4da66d4e,
        64'h8afd13cf8e6fb054, 64'hf5e1c9011d5ed849, 64'he34e091c5126c8af, 64'had67ee7530a398f6,
        64'h43b24dec2e82c75a, 64'h75da99c1287cd48d, 64'h92e81cdb3783f689, 64'ha3dd217cc537cecd,
        64'h60543c50de970553, 64'h93f73f54aaf2426a, 64'ha91b62737e7a725d, 64'hf19d4507538732e2,
        64'h77e4dfc20f9ea156, 64'h7d229ccdb4d31dc6, 64'h1b346a98037f87e5, 64'hedf4c615a4b29e94,
        64'h4093286094110662, 64'hb0114ee85ae78063, 64'h6ff1d0d6b672e78b, 64'h6dcf96d591909250,
        64'hdfe09e3eec9567e8, 64'h3214582b4827f97c, 64'hb46dc2ee143e6ac8, 64'hf6c0ac8da7cd1971,
        64'hebb60c10cd8901e4, 64'hf7df8f023abcad92, 64'h9c52d3d2c217a0b2, 64'h6b8d5cd0f8ab0d20,
        64'h3777f7a29b8fa734, 64'h011f238f9d71b4e3, 64'hc1b75b2f3c42be45, 64'h5de588fdfe551ef7,
        64'h6eeef3592b035368, 64'haa3a07ffc4e9b365, 64'hecebe59a39c32a77, 64'h5ba742f8976e8187,
        64'h4b4a48e0b22d0e11, 64'hddded83dcb771233, 64'ha59feb79ac0c51bd, 64'hc7f5912a55792135
        };
logic [0:255][63:0] T5 = {64'h6d6ae04668a9b08a, 64'h3ab3f04b0be8c743, 64'he51e166b54b3c908, 64'hbe90a9eb35c2f139,
        64'hb2c7066637f2bec1, 64'haa6945613392202c, 64'h9a28c36f3b5201eb, 64'hddce5a93ab536994,
        64'h0e34133ef6382827, 64'h52a02ba1ec55048b, 64'ha2f88f97c4b2a177, 64'h8640e513ca2251a5,
        64'hcdf1d36258137622, 64'hfe6cb708dedf8ddb, 64'h8a174a9ec8121e5d, 64'h679896036b81560e,
        64'h59ed033395795fee, 64'h1dd778ab8b74edaf, 64'hee533ef92d9f926d, 64'h2a8c79baf8a8d8f5,
        64'h6bcf398e69b119f6, 64'he20491742fafdd95, 64'h276488e0809c2aec, 64'hea955b82d88f5cce,
        64'h7102c63a99d9e0c4, 64'hf9763017a5c39946, 64'h429fa2501f151b3d, 64'h4659c72bea05d59e,
        64'h984b7fdccf5a6634, 64'hf742232953fbb161, 64'h3041860e08c021c7, 64'h747bfd9616cd9386,
        64'h4bb1367192312787, 64'h1b72a1638a6c44d3, 64'h4a0e68a6e8359a66, 64'h169a5039f258b6ca,
        64'hb98a2ef44edee5a4, 64'hd9083fe85e43a737, 64'h967f6ce239624e13, 64'h8874f62d3c1a7982,
        64'h3c1629830af06e3f, 64'h9165ebfd427e5a8e, 64'hb5dd81794ceeaa5c, 64'h0de8f15a7834f219,
        64'h70bd98ede3dd5d25, 64'haccc9ca9328a8950, 64'h56664eda1945ca28, 64'h221db34c0f8859ae,
        64'h26dbd637fa98970d, 64'h1acdffb4f068f932, 64'h4585254f64090fa0, 64'h72de245e17d53afa,
        64'h1546b25d7c546cf4, 64'h207e0ffffb803e71, 64'hfaaad2732bcf4378, 64'hb462dfae36ea17bd,
        64'hcf926fd1ac1b11fd, 64'he0672dc7dba7ba4a, 64'hd3fa49ad5d6b41b3, 64'h8ba81449b216a3bc,
        64'h14f9ec8a0650d115, 64'h40fc1ee3eb1d7ce2, 64'h23a2ed9b758ce44f, 64'h782c521b14fddc7e,
        64'h1c68267cf170504e, 64'hbcf31558c1ca96e6, 64'ha781b43b4ba6d235, 64'hf6fd7dfe29ff0c80,
        64'hb0a4bad5c3fad91e, 64'hd199f51ea963266c, 64'h414340349119c103, 64'h5405f269ed4dadf7,
        64'habd61bb649969dcd, 64'h6813dbeae7bdc3c8, 64'h65fb2ab09f8931d1, 64'hf1e7fae152e3181d,
        64'hc1a67cef5a2339da, 64'h7a4feea8e0f5bba1, 64'h1e0b9acf05783791, 64'h5b8ebf8061713831,
        64'h80e53cdbcb3af8d9, 64'h7e898bd315e57502, 64'hc6bcfbf0213f2d47, 64'h95a38e86b76e942d,
        64'h092e94218d243cba, 64'h8339debf453622e7, 64'hb11be402b9fe64ff, 64'h57d9100d634177c9,
        64'hcc4e8db52217cbc3, 64'h3b0cae9c71ec7aa2, 64'hfb158ca451cbfe99, 64'h2b33276d82ac6514,
        64'h01bf5ed77a04bde1, 64'hc5601994af33f779, 64'h75c4a3416cc92e67, 64'hf3844652a6eb7fc2,
        64'h3487e375fdd0ef64, 64'h18ae430704609eed, 64'h4d14efb993298efb, 64'h815a620cb13e4538,
        64'h125c354207487869, 64'h9eeea614ce42cf48, 64'hce2d3106d61fac1c, 64'hbbe99247bad6827b,
        64'h071a871f7b1c149d, 64'h2e4a1cc10db81656, 64'h77a71ff298c149b8, 64'h06a5d9c80118a97c,
        64'had73c27e488e34b1, 64'h443a7b981e0db241, 64'he3bbcfa355ab6074, 64'h0af276450328e684,
        64'h73617a896dd1871b, 64'h58525de4ef7de20f, 64'hb7be3dcab8e6cd83, 64'h19111dd07e64230c,
        64'h842359a03e2a367a, 64'h103f89f1f3401fb6, 64'hdc710444d157d475, 64'hb835702334da5845,
        64'h4320fc876511a6dc, 64'hd026abc9d3679b8d, 64'h17250eee885c0b2b, 64'h90dab52a387ae76f,
        64'h31fed8d972c49c26, 64'h89cba8fa461ec463, 64'h2ff5421677bcabb7, 64'h396f122f85e41d7d,
        64'ha09b332430bac6a8, 64'hc888e8ced7070560, 64'haeaf201ac682ee8f, 64'h1180d7268944a257,
        64'hf058a43628e7a5fc, 64'hbd4c4b8fbbce2b07, 64'ha1246df34abe7b49, 64'h7d5569b79be9af3c,
        64'ha9b5a705bd9efa12, 64'hdb6b835baa4bc0e8, 64'h05793bac8f147342, 64'h21c1512881848390,
        64'hfdb0556c50d357e5, 64'h613d4fcb6a99ff72, 64'h03dce2648e0cda3e, 64'he949b9e6568386f0,
        64'hfc0f0bbb2ad7ea04, 64'h6a70675913b5a417, 64'h7f36d5046fe1c8e3, 64'h0c57af8d02304ff8,
        64'h32223abdfcc84618, 64'h0891caf6f720815b, 64'ha63eeaec31a26fd4, 64'h2507345374944d33,
        64'h49d28ac266394058, 64'hf5219f9aa7f3d6be, 64'h2d96fea583b4cc68, 64'h5a31e1571b7585d0,
        64'h8ed12fe53d02d0fe, 64'hdfade6205f5b0e4b, 64'h4cabb16ee92d331a, 64'h04c6657bf510cea3,
        64'hd73c2cd6a87b8f10, 64'he1d87310a1a307ab, 64'h6cd5be9112ad0d6b, 64'h97c032354366f3f2,
        64'hd4e0ceb22677552e, 64'h0000000000000000, 64'h29509bde76a402cb, 64'hc27a9e8bd42fe3e4,
        64'h5ef7842cee654b73, 64'haf107ecdbc86536e, 64'h3fcacbe784fcb401, 64'hd55f90655c73e8cf,
        64'he6c2f40fdabf1336, 64'he8f6e7312c873b11, 64'heb2a0555a28be12f, 64'he4a148bc2eb774e9,
        64'h9b979db84156bc0a, 64'h6eb60222e6a56ab4, 64'h87ffbbc4b026ec44, 64'hc703a5275b3b90a6,
        64'h47e699fc9001687f, 64'h9c8d1aa73a4aa897, 64'h7cea3760e1ed12dd, 64'h4ec80ddd1d2554c5,
        64'h13e36b957d4cc588, 64'h5d2b66486069914d, 64'h92b90999cc7280b0, 64'h517cc9c56259deb5,
        64'hc937b619ad03b881, 64'hec30824ad997f5b2, 64'ha45d565fc5aa080b, 64'hd6837201d27f32f1,
        64'h635ef3789e9198ad, 64'h531f75769651b96a, 64'h4f77530a6721e924, 64'h486dd4151c3dfdb9,
        64'h5f48dafb9461f692, 64'h375b011173dc355a, 64'h3da9775470f4d3de, 64'h8d0dcd81b30e0ac0,
        64'h36e45fc609d888bb, 64'h55baacbe97491016, 64'h8cb29356c90ab721, 64'h76184125e2c5f459,
        64'h99f4210bb55edbd5, 64'h6f095cf59ca1d755, 64'h9f51f8c3b44672a9, 64'h3538bda287d45285,
        64'h50c39712185d6354, 64'hf23b1885dcefc223, 64'h79930ccc6ef9619f, 64'hed8fdc9da3934853,
        64'hcb540aaa590bdf5e, 64'h5c94389f1a6d2cac, 64'he77daad8a0bbaed7, 64'h28efc5090ca0bf2a,
        64'hbf2ff73c4fc64cd8, 64'hb37858b14df60320, 64'hf8c96ec0dfc724a7, 64'h828680683f329f06,
        64'h941cd051cd6a29cc, 64'hc3c5c05cae2b5e05, 64'hb601631dc2e27062, 64'hc01922382027843b,
        64'h24b86a840e90f0d2, 64'hd245177a276ffc52, 64'h0f8b4de98c3c95c6, 64'h3e759530fef809e0,
        64'h0b4d2892792c5b65, 64'hc4df4743d5374a98, 64'ha5e20888bfaeb5ea, 64'hba56cc90c0d23f9a,
        64'h38d04cf8ffe0a09c, 64'h62e1adafe495254c, 64'h0263bcb3f40867df, 64'hcaeb547d230f62bf,
        64'h6082111c109d4293, 64'hdad4dd8cd04f7d09, 64'hefec602e579b2f8c, 64'h1fb4c4187f7c8a70,
        64'hffd3e9dfa4db303a, 64'h7bf0b07f9af10640, 64'hf49ec14dddf76b5f, 64'h8f6e713247066d1f,
        64'h339d646a86ccfbf9, 64'h64447467e58d8c30, 64'h2c29a072f9b07189, 64'hd8b7613f24471ad6,
        64'h6627c8d41185ebef, 64'ha347d140beb61c96, 64'hde12b8f7255fb3aa, 64'h9d324470404e1576,
        64'h9306574eb6763d51, 64'ha80af9d2c79a47f3, 64'h859c0777442e8b9b, 64'h69ac853d9db97e29
        };
        logic [0:255][63:0] T6 = {64'hc3407dfc2de6377e, 64'h5b9e93eea4256f77, 64'hadb58fdd50c845e0, 64'h5219ff11a75bed86,
        64'h356b61cfd90b1de9, 64'hfb8f406e25abe037, 64'h7a5a0231c0f60796, 64'h9d3cd216e1f5020b,
        64'h0c6550fb6b48d8f3, 64'hf57508c427ff1c62, 64'h4ad35ffa71cb407d, 64'h6290a2da1666aa6d,
        64'he284ec2349355f9f, 64'hb3c307c53d7c84ec, 64'h05e23c0468365a02, 64'h190bac4d6c9ebfa8,
        64'h94bbbee9e28b80fa, 64'ha34fc777529cb9b5, 64'hcc7b39f095bcd978, 64'h2426addb0ce532e3,
        64'h7e79329312ce4fc7, 64'hab09a72eebec2917, 64'hf8d15499f6b9d6c2, 64'h1a55b8babf8c895d,
        64'hdb8add17fb769a85, 64'hb57f2f368658e81b, 64'h8acd36f18f3f41f6, 64'h5ce3b7bba50f11d3,
        64'h114dcc14d5ee2f0a, 64'hb91a7fcded1030e8, 64'h81d5425fe55de7a1, 64'hb6213bc1554adeee,
        64'h80144ef95f53f5f2, 64'h1e7688186db4c10c, 64'h3b912965db5fe1bc, 64'hc281715a97e8252d,
        64'h54a5d7e21c7f8171, 64'h4b12535ccbc5522e, 64'h1d289cefbea6f7f9, 64'h6ef5f2217d2e729e,
        64'he6a7dc819b0d17ce, 64'h1b94b41c05829b0e, 64'h33d7493c622f711e, 64'hdcf7f942fa5ce421,
        64'h600fba8b7f7a8ecb, 64'h46b60f011a83988e, 64'h235b898e0dcf4c47, 64'h957ab24f588592a9,
        64'h4354330572b5c28c, 64'ha5f3ef84e9b8d542, 64'h8c711e02341b2d01, 64'h0b1874ae6a62a657,  
        64'h1213d8e306fc19ff, 64'hfe6d7c6a4d9dba35, 64'h65ed868f174cd4c9, 64'h88522ea0e6236550,
        64'h899322065c2d7703, 64'hc01e690bfef4018b, 64'h915982ed8abddaf8, 64'hbe675b98ec3a4e4c,
        64'ha996bf7f82f00db1, 64'he1daf8d49a27696a, 64'h2effd5d3dc8986e7, 64'hd153a51f2b1a2e81,
        64'h18caa0ebd690adfb, 64'h390e3134b243c51a, 64'h2778b92cdff70416, 64'h029f1851691c24a6,
        64'h5e7cafeacc133575, 64'hfa4e4cc89fa5f264, 64'h5a5f9f481e2b7d24, 64'h484c47ab18d764db,
        64'h400a27f2a1a7f479, 64'haeeb9b2a83da7315, 64'h721c626879869734, 64'h042330a2d2384851,
        64'h85f672fd3765aff0, 64'hba446b3a3e02061d, 64'h73dd6ecec3888567, 64'hffac70ccf793a866,
        64'hdfa9edb5294ed2d4, 64'h6c6aea7014325638, 64'h834a5a0e8c41c307, 64'hcdba35562fb2cb2b,
        64'h0ad97808d06cb404, 64'h0f3b440cb85aee06, 64'he5f9c876481f213b, 64'h98deee1289c35809,
        64'h59018bbfcd394bd1, 64'he01bf47220297b39, 64'hde68e1139340c087, 64'h9fa3ca4788e926ad,
        64'hbb85679c840c144e, 64'h53d8f3b71d55ffd5, 64'h0da45c5dd146caa0, 64'h6f34fe87c72060cd,
        64'h57fbc315cf6db784, 64'hcee421a1fca0fdde, 64'h3d2d0196607b8d4b, 64'h642c8a29ad42c69a,
        64'h14aff010bdd87508, 64'hac74837beac657b3, 64'h3216459ad821634d, 64'h3fb219c70967a9ed,
        64'h06bc28f3bb246cf7, 64'hf2082c9126d562c6, 64'h66b39278c45ee23c, 64'hbd394f6f3f2878b9,
        64'hfd33689d9e8f8cc0, 64'h37f4799eb017394f, 64'h108cc0b26fe03d59, 64'hda4bd1b1417888d6,
        64'hb09d1332ee6eb219, 64'h2f3ed975668794b4, 64'h58c0871977375982, 64'h7561463d78ace990,
        64'h09876cff037e82f1, 64'h7fb83e35a8c05d94, 64'h26b9b58a65f91645, 64'hef20b07e9873953f,
        64'h3148516d0b3355b8, 64'h41cb2b541ba9e62a, 64'h790416c613e43163, 64'ha011d380818e8f40,
        64'h3a5025c36151f3ef, 64'hd57095bdf92266d0, 64'h498d4b0da2d97688, 64'h8b0c3a57353153a5,
        64'h21c491df64d368e1, 64'h8f2f0af5e7091bf4, 64'h2da1c1240f9bb012, 64'hc43d59a92ccc49da,
        64'hbfa6573e56345c1f, 64'h828b56a8364fd154, 64'h9a41f643e0df7caf, 64'hbcf843c985266aea,
        64'h2b1de9d7b4bfdce5, 64'h20059d79dedd7ab2, 64'h6dabe6d6ae3c446b, 64'h45e81bf6c991ae7b,
        64'h6351ae7cac68b83e, 64'ha432e32253b6c711, 64'hd092a9b991143cd2, 64'hcac711032e98b58f,
        64'hd8d4c9e02864ac70, 64'hc5fc550f96c25b89, 64'hd7ef8dec903e4276, 64'h67729ede7e50f06f,
        64'heac28c7af045cf3d, 64'hb15c1f945460a04a, 64'h9cfddeb05bfb1058, 64'h93c69abce3a1fe5e,
        64'heb0380dc4a4bdd6e, 64'hd20db1e8f8081874, 64'h229a8528b7c15e14, 64'h44291750739fbc28,
        64'hd3ccbd4e42060a27, 64'hf62b1c33f4ed2a97, 64'h86a8660ae4779905, 64'hd62e814a2a305025,
        64'h477703a7a08d8add, 64'h7b9b0e977af815c5, 64'h78c51a60a9ea2330, 64'ha6adfb733aaae3b7,
        64'h97e5aa1e3199b60f, 64'h0000000000000000, 64'hf4b404629df10e31, 64'h5564db44a6719322,
        64'h9207961a59afec0d, 64'h9624a6b88b97a45c, 64'h363575380a192b1c, 64'h2c60cd82b595a241,
        64'h7d272664c1dc7932, 64'h7142769faa94a1c1, 64'ha1d0df263b809d13, 64'h1630e841d4c451ae,
        64'hc1df65ad44fa13d8, 64'h13d2d445bcf20bac, 64'hd915c546926abe23, 64'h38cf3d92084dd749,
        64'he766d0272103059d, 64'hc7634d5effde7f2f, 64'h077d2455012a7ea4, 64'hedbfa82ff16fb199,
        64'haf2a978c39d46146, 64'h42953fa3c8bbd0df, 64'hcb061da59496a7dc, 64'h25e7a17db6eb20b0,
        64'h34aa6d6963050fba, 64'ha76cf7d580a4f1e4, 64'hf7ea10954ee338c4, 64'hfcf2643b24819e93,
        64'hcf252d0746aeef8d, 64'h4ef06f58a3f3082c, 64'h563acfb37563a5d7, 64'h5086e740ce47c920,
        64'h2982f186dda3f843, 64'h87696aac5e798b56, 64'h5d22bb1d1f010380, 64'h035e14f7d31236f5,
        64'h3cec0d30da759f18, 64'hf3c920379cdb7095, 64'hb8db736b571e22bb, 64'hdd36f5e44052f672,
        64'haac8ab8851e23b44, 64'ha857b3d938fe1fe2, 64'h17f1e4e76eca43fd, 64'hec7ea4894b61a3ca,
        64'h9e62c6e132e734fe, 64'hd4b1991b432c7483, 64'h6ad6c283af163acf, 64'h1ce9904904a8e5aa,
        64'h5fbda34c761d2726, 64'hf910583f4cb7c491, 64'hc6a241f845d06d7c, 64'h4f3163fe19fd1a7f,
        64'he99c988d2357f9c8, 64'h8eee06535d0709a7, 64'h0efa48aa0254fc55, 64'hb4be23903c56fa48,
        64'h763f52caabbedf65, 64'heee1bcd8227d876c, 64'he345e085f33b4dcc, 64'h3e731561b369bbbe,
        64'h2843fd2067adea10, 64'h2adce5710eb1ceb6, 64'hb7e03767ef44ccbd, 64'h8db012a48e153f52,
        64'h61ceb62dc5749c98, 64'he85d942b9959eb9b, 64'h4c6f7709caef2c8a, 64'h84377e5b8d6bbda3,
        64'h30895dcbb13d47eb, 64'h74a04a9bc2a2fbc3, 64'h6b17ce251518289c, 64'he438c4d0f2113368,
        64'h1fb784bed7bad35f, 64'h9b80fae55ad16efc, 64'h77fe5e6c11b0cd36, 64'hc858095247849129,
        64'h08466059b97090a2, 64'h01c10ca6ba0e1253, 64'h6988d6747c040c3a, 64'h6849dad2c60a1e69,
        64'h5147ebe67449db73, 64'hc99905f4fd8a837a, 64'h991fe2b433cd4a5a, 64'hf09734c04fc94660,
        64'ha28ecbd1e892abe6, 64'hf1563866f5c75433, 64'h4dae7baf70e13ed9, 64'h7ce62ac27bd26b61,
        64'h70837a39109ab392, 64'h90988e4b30b3c8ab, 64'hb2020b63877296bf, 64'h156efcb607d6675b
        };
logic [0:255][63:0] T7 = {64'he63f55ce97c331d0, 64'h25b506b0015bba16, 64'hc8706e29e6ad9ba8, 64'h5b43d3775d521f6a,
        64'h0bfa3d577035106e, 64'hab95fc172afb0e66, 64'hf64b63979e7a3276, 64'hf58b4562649dad4b,
        64'h48f7c3dbae0c83f1, 64'hff31916642f5c8c5, 64'hcbb048dc1c4a0495, 64'h66b8f83cdf622989,
        64'h35c130e908e2b9b0, 64'h7c761a61f0b34fa1, 64'h3601161cf205268d, 64'h9e54ccfe2219b7d6,
        64'h8b7d90a538940837, 64'h9cd403588ea35d0b, 64'hbc3c6fea9ccc5b5a, 64'he5ff733b6d24aeed,
        64'hceed22de0f7eb8d2, 64'hec8581cab1ab545e, 64'hb96105e88ff8e71d, 64'h8ca03501871a5ead,
        64'h76ccce65d6db2a2f, 64'h5883f582a7b58057, 64'h3f7be4ed2e8adc3e, 64'h0fe7be06355cd9c9,
        64'hee054e6c1d11be83, 64'h1074365909b903a6, 64'h5dde9f80b4813c10, 64'h4a770c7d02b6692c,
        64'h5379c8d5d7809039, 64'hb4067448161ed409, 64'h5f5e5026183bd6cd, 64'he898029bf4c29df9,
        64'h7fb63c940a54d09c, 64'hc5171f897f4ba8bc, 64'ha6f28db7b31d3d72, 64'h2e4f3be7716eaa78,
        64'h0d6771a099e63314, 64'h82076254e41bf284, 64'h2f0fd2b42733df98, 64'h5c9e76d3e2dc49f0,
        64'h7aeb569619606cdb, 64'h83478b07b2468764, 64'hcfadcb8d5923cd32, 64'h85dac7f05b95a41e,
        64'hb5469d1b4043a1e9, 64'hb821ecbbd9a592fd, 64'h1b8e0b0e798c13c8, 64'h62a57b6d9a0be02e,
        64'hfcf1b793b81257f8, 64'h9d94ea0bd8fe28eb, 64'h4cea408aeb654a56, 64'h23284a47e888996c,
        64'h2d8f1d128b893545, 64'hf4cbac3132c0d8ab, 64'hbd7c86b9ca912eba, 64'h3a268eef3dbe6079,
        64'hf0d62f6077a9110c, 64'h2735c916ade150cb, 64'h89fd5f03942ee2ea, 64'h1acee25d2fd16628,
        64'h90f39bab41181bff, 64'h430dfe8cde39939f, 64'hf70b8ac4c8274796, 64'h1c53aeaac6024552,
        64'h13b410acf35e9c9b, 64'ha532ab4249faa24f, 64'h2b1251e5625a163f, 64'hd7e3e676da4841c7,
        64'ha7b264e4e5404892, 64'hda8497d643ae72d3, 64'h861ae105a1723b23, 64'h38a6414991048aa4,
        64'h6578dec92585b6b4, 64'h0280cfa6acbaeadd, 64'h88bdb650c273970a, 64'h9333bd5ebbff84c2,
        64'h4e6a8f2c47dfa08b, 64'h321c954db76cef2a, 64'h418d312a72837942, 64'hb29b38bfffcdf773,
        64'h6c022c38f90a4c07, 64'h5a033a240b0f6a8a, 64'h1f93885f3ce5da6f, 64'hc38a537e96988bc6,
        64'h39e6a81ac759ff44, 64'h29929e43cee0fce2, 64'h40cdd87924de0ca2, 64'he9d8ebc8a29fe819,
        64'h0c2798f3cfbb46f4, 64'h55e484223e53b343, 64'h4650948ecd0d2fd8, 64'h20e86cb2126f0651,
        64'h6d42c56baf5739e7, 64'ha06fc1405ace1e08, 64'h7babbfc54f3d193b, 64'h424d17df8864e67f,
        64'hd8045870ef14980e, 64'hc6d7397c85ac3781, 64'h21a885e1443273b1, 64'h67f8116f893f5c69,
        64'h24f5efe35706cff6, 64'hd56329d076f2ab1a, 64'h5e1eb9754e66a32d, 64'h28d2771098bd8902,
        64'h8f6013f47dfdc190, 64'h17a993fdb637553c, 64'he0a219397e1012aa, 64'h786b9930b5da8606,
        64'h6e82e39e55b0a6da, 64'h875a0856f72f4ec3, 64'h3741ff4fa458536d, 64'hac4859b3957558fc,
        64'h7ef6d5c75c09a57c, 64'hc04a758b6c7f14fb, 64'hf9acdd91ab26ebbf, 64'h7391a467c5ef9668,
        64'h335c7c1ee1319aca, 64'ha91533b18641e4bb, 64'he4bf9a683b79db0d, 64'h8e20faa72ba0b470,
        64'h51f907737b3a7ae4, 64'h2268a314bed5ec8c, 64'hd944b123b949edee, 64'h31dcb3b84d8b7017,
        64'hd3fe65279f218860, 64'h097af2f1dc8ffab3, 64'h9b09a6fc312d0b91, 64'hcc6ded78a3c4520f,
        64'h3481d9ba5ebfcc50, 64'h4f2a667f1182d56b, 64'hdfd9fdd4509ace94, 64'h26752045fbbc252b,
        64'hbffc491f662bc467, 64'hdd593272fc202449, 64'h3cbbc218d46d4303, 64'h91b372f817456e1f,
        64'h681faf69bc6385a0, 64'hb686bbeebaa43ed4, 64'h1469b5084cd0ca01, 64'h98c98009cbca94ac,
        64'h6438379a73d8c354, 64'hc2caba2dc0c5fe26, 64'h3e3b0dbe78d7a9de, 64'h50b9ee202d670f04,
        64'h4590b27b37eab0e5, 64'h6025b4cb36b10af3, 64'hfb2c1237079c0162, 64'ha12f28130c936be8,
        64'h4b37e52e54eb1ccc, 64'h083a1ba28ad28f53, 64'hc10a9cd83a22611b, 64'h9f1425ad7444c236,
        64'h069d4cf7e9d3237a, 64'hedc56899e7f621be, 64'h778c273680865fcf, 64'h309c5aeb1bd605f7,
        64'h8de0dc52d1472b4d, 64'hf8ec34c2fd7b9e5f, 64'hea18cd3d58787724, 64'haad515447ca67b86,
        64'h9989695a9d97e14c, 64'h0000000000000000, 64'hf196c63321f464ec, 64'h71116bc169557cb5,
        64'haf887f466f92c7c1, 64'h972e3e0ffe964d65, 64'h190ec4a8d536f915, 64'h95aef1a9522ca7b8,
        64'hdc19db21aa7d51a9, 64'h94ee18fa0471d258, 64'h8087adf248a11859, 64'hc457f6da2916dd5c,
        64'hfa6cfb6451c17482, 64'hf256e0c6db13fbd1, 64'h6a9f60cf10d96f7d, 64'h4daaa9d9bd383fb6,
        64'h03c026f5fae79f3d, 64'hde99148706c7bb74, 64'h2a52b8b6340763df, 64'h6fc20acd03edd33a,
        64'hd423c08320afdefa, 64'hbbe1ca4e23420dc0, 64'h966ed75ca8cb3885, 64'heb58246e0e2502c4,
        64'h055d6a021334bc47, 64'ha47242111fa7d7af, 64'he3623fcc84f78d97, 64'h81c744a11efc6db9,
        64'haec8961539cfb221, 64'hf31609958d4e8e31, 64'h63e5923ecc5695ce, 64'h47107ddd9b505a38,
        64'ha3afe7b5a0298135, 64'h792b7063e387f3e6, 64'h0140e953565d75e0, 64'h12f4f9ffa503e97b,
        64'h750ce8902c3cb512, 64'hdbc47e8515f30733, 64'h1ed3610c6ab8af8f, 64'h5239218681dde5d9,
        64'he222d69fd2aaf877, 64'hfe71783514a8bd25, 64'hcaf0a18f4a177175, 64'h61655d9860ec7f13,
        64'he77fbc9dc19e4430, 64'h2ccff441ddd440a5, 64'h16e97aaee06a20dc, 64'ha855dae2d01c915b,
        64'h1d1347f9905f30b2, 64'hb7c652bdecf94b34, 64'hd03e43d265c6175d, 64'hfdb15ec0ee4f2218,
        64'h57644b8492e9599e, 64'h07dda5a4bf8e569a, 64'h54a46d71680ec6a3, 64'h5624a2d7c4b42c7e,
        64'hbebca04c3076b187, 64'h7d36f332a6ee3a41, 64'h3b6667bc6be31599, 64'h695f463aea3ef040,
        64'had08b0e0c3282d1c, 64'hb15b1e4a052a684e, 64'h44d05b2861b7c505, 64'h15295c5b1a8dbfe1,
        64'h744c01c37a61c0f2, 64'h59c31cd1f1e8f5b7, 64'hef45a73f4b4ccb63, 64'h6bdf899c46841a9d,
        64'h3dfb2b4b823036e3, 64'ha2ef0ee6f674f4d5, 64'h184e2dfb836b8cf5, 64'h1134df0a5fe47646,
        64'hbaa1231d751f7820, 64'hd17eaa81339b62bd, 64'hb01bf71953771dae, 64'h849a2ea30dc8d1fe,
        64'h705182923f080955, 64'h0ea757556301ac29, 64'h041d83514569c9a7, 64'h0abad4042668658e,
        64'h49b72a88f851f611, 64'h8a3d79f66ec97dd7, 64'hcd2d042bf59927ef, 64'hc930877ab0f0ee48,
        64'h9273540deda2f122, 64'hc797d02fd3f14261, 64'he1e2f06a284d674a, 64'hd2be8c74c97cfd80,
        64'h9a494faf67707e71, 64'hb3dbd1eca9908293, 64'h72d14d3493b2e388, 64'hd6a30f258c153427
};
 

always @(posedge clk_i or negedge rstn_i)
if(!rstn_i)
  begin
   valid_o <= '0;   
  end
else 
  begin     
   valid_o <= valid_i;
  end 
 always_comb
    begin
    internal[0] = T0[(state[0])]  ^ T1[(state[8])] ^ T2[(state[16])] ^ T3[(state[24])] ^
            T4[(state[32])] ^ T5[(state[40])] ^ T6[(state[48])] ^ T7[(state[56])];
    internal[1] = T0[(state[1])] ^ T1[(state[9])] ^ T2[(state[17])] ^ T3[(state[25])] ^
            T4[(state[33])] ^ T5[(state[41])] ^ T6[(state[49])] ^ T7[(state[57])];
    internal[2] = T0[(state[2])] ^ T1[(state[10])] ^ T2[(state[18])] ^ T3[(state[26])] ^
            T4[(state[34])] ^ T5[(state[42])] ^ T6[(state[50])] ^ T7[(state[58])];
    internal[3] = T0[(state[3])] ^ T1[(state[11])] ^ T2[(state[19])] ^ T3[(state[27])] ^
            T4[(state[35])] ^ T5[(state[43])] ^ T6[(state[51])] ^ T7[(state[59])];
    internal[4] = T0[(state[4])] ^ T1[(state[12])] ^ T2[(state[20])] ^ T3[(state[28])] ^
            T4[(state[36])] ^ T5[(state[44])] ^ T6[(state[52])] ^ T7[(state[60])];
    internal[5] = T0[(state[5])] ^ T1[(state[13])] ^ T2[(state[21])] ^ T3[(state[29])] ^
            T4[(state[37])] ^ T5[(state[45])] ^ T6[(state[53])] ^ T7[(state[61])];
    internal[6] = T0[(state[6])] ^ T1[(state[14])] ^ T2[(state[22])] ^ T3[(state[30])] ^
            T4[(state[38])] ^ T5[(state[46])] ^ T6[(state[54])] ^ T7[(state[62])];
    internal[7] = T0[(state[7])] ^ T1[(state[15])] ^ T2[(state[23])] ^ T3[(state[31])] ^
            T4[(state[39])] ^ T5[(state[47])] ^ T6[(state[55])] ^ T7[(state[63])];
     end
assign state_f = lps_n_i ^ lps_m_i;

always_comb
for(int i = 0; i < 64 ; i++)
   state[i] <= state_f[8*i+7-:8];

always @(posedge clk_i or negedge rstn_i)
if(!rstn_i)
  lps_o   <= '0;                
else if(valid_i)
       lps_o <= {internal[7],internal[6],internal[5],internal[4],internal[3],internal[2],internal[1],internal[0]};

endmodule